/*
 * Módulo: ula_8bits
 * Função: ULA que realiza 8 operações em paralelo e seleciona uma saída.
 */
module ula_8bits (
    input [7:0] a,
    input [7:0] b,
    input [2:0] sel_op,
    output [7:0] resultado_ula
    // Adicione aqui as saídas para os flags (Zero, Overflow, etc.)
);
    // Fios para guardar o resultado de CADA operação
    wire [7:0] res_soma, res_sub, res_mult, res_div;
    wire [7:0] res_and, res_or, res_xor, res_not;

    // --- 1. INSTANCIE SEUS MÓDULOS DE OPERAÇÃO ---
    // Eles estão todos trabalhando em paralelo, o tempo todo.
    // **IMPORTANTE: Ajuste os nomes dos módulos e das portas (.a, .b, .soma, etc.)
    // para corresponderem exatamente aos que você criou!**

    somadorde8bits      MOD_SOMA (.A(a), .B(b), .S(res_soma));
    subtrator_8bits    MOD_SUB  (.A(a), .B(b), .S(res_sub));
    multiplicador_8bits MOD_MULT (.a(a), .b(b), .s(res_mult)); // Módulo sequencial que você fará
    divisor_8bits      MOD_DIV  (.a(a), .b(b), .s(res_div));   // Módulo sequencial que você fará
    opLogicoAND          MOD_AND  (.A(a), .B(b), .S(res_and));
    opLogicoOR           MOD_OR   (.A(a), .B(b), .S(res_or));
    opLogicoXOR          MOD_XOR  (.A(a), .B(b), .S(res_xor));
    opLogicoNOT          MOD_NOT  (.A(a), .S(res_not)); // NOT só precisa de uma entrada

    // --- 2. INSTANCIE O MUX SELETOR ---
    // O MUX seleciona qual dos resultados vai para a saída final.
    mux_8para1_8bits MUX_SELETOR (
        .in0(res_soma),
        .in1(res_sub),
        .in2(res_mult),
        .in3(res_div),
        .in4(res_and),
        .in5(res_or),
        .in6(res_xor),
        .in7(res_not),
        .sel(sel_op),
        .out(resultado_ula)
    );

endmodule
